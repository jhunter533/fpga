module linear_layer #(
  parameter INPUT=x,
  parameter OUTPUT=y,
)(
  input clk,
  imput rsk,
  input ...
  output ...
);
  localparam TOTAL_WIDTH=16;

